// Broderick Bownds
// brbownds@hmc.edu
// 9/6/2025

module lab2_bb( input  logic reset,
				input  logic [3:0] s0,
				input  logic [3:0] s1,
				output logic [5:0] led,
				output logic [6:0] seg);	

	
	endmodule